module main
import cli


fn main() {
	cli.start_cli()
}
