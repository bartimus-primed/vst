module implant

// detect os

// start beacon

// wait for tasks
