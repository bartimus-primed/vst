module c2

import os

// detect os

pub fn get_os() string {
	return os.user_os()
}


// start listener

// interact

// schedule tasks