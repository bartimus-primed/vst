module main

import c2

fn main() {
	println(c2.get_os())
}