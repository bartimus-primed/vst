module linux