module cli

import c2

pub fn start_cli() {
	c2.start_c2()
}